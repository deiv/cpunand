
Library IEEE;
USE IEEE.Std_logic_1164.all;

entity DFF is
   port(
      q   : out std_logic;
      clk : in std_logic;
      d   : in std_logic
   );
end DFF;

architecture Behavioral of DFF is
begin
 process(clk)
 begin
    if(rising_edge(clk)) then
        q <= d;
    end if;
 end process;
end Behavioral;


Library IEEE;
USE IEEE.Std_logic_1164.all;

entity register1 is port(
    d   : in std_logic;
    ld  : in std_logic; -- load/enable.
    clk : in std_logic; -- clock.
    q   : out std_logic -- output.
);
end register1;

architecture description of register1 IS

begin
    process(clk)
    begin
        if rising_edge(clk) then
            if ld = '1' then
                q <= d;
            end if;
        end if;
    end process;
end description;


library ieee;
use ieee.std_logic_1164.all;

entity register32 is port(
    d   : in std_logic_vector(31 downto 0);
    ld  : in std_logic;                     -- load/enable.
    clk : in std_logic;                     -- clock.
    q   : out std_logic_vector(31 downto 0) -- output
);
end register32;

architecture description of register32 is

begin
    process(clk)
    begin
        if rising_edge(clk) then
            if ld = '1' then
                q <= d;
            end if;
        end if;
    end process;
end description;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;

-- A 128x8 single-port RAM in VHDL
entity Single_port_RAM_VHDL is
port(
 RAM_ADDR: in std_logic_vector(6 downto 0); -- Address to write/read RAM
 RAM_DATA_IN: in std_logic_vector(7 downto 0); -- Data to write into RAM
 RAM_WR: in std_logic; -- Write enable
 RAM_CLOCK: in std_logic; -- clock input for RAM
 RAM_DATA_OUT: out std_logic_vector(7 downto 0) -- Data output of RAM
);
end Single_port_RAM_VHDL;

architecture Behavioral of Single_port_RAM_VHDL is
-- define the new type for the 128x8 RAM
type RAM_ARRAY is array (0 to 127 ) of std_logic_vector (7 downto 0);
-- initial values in the RAM
signal RAM: RAM_ARRAY :=(
   x"55",x"66",x"77",x"67",-- 0x00:
   x"99",x"00",x"00",x"11",-- 0x04:
   x"00",x"00",x"00",x"00",-- 0x08:
   x"00",x"00",x"00",x"00",-- 0x0C:
   x"00",x"00",x"00",x"00",-- 0x10:
   x"00",x"00",x"00",x"00",-- 0x14:
   x"00",x"00",x"00",x"00",-- 0x18:
   x"00",x"00",x"00",x"00",-- 0x1C:
   x"00",x"00",x"00",x"00",-- 0x20:
   x"00",x"00",x"00",x"00",-- 0x24:
   x"00",x"00",x"00",x"00",-- 0x28:
   x"00",x"00",x"00",x"00",-- 0x2C:
   x"00",x"00",x"00",x"00",-- 0x30:
   x"00",x"00",x"00",x"00",-- 0x34:
   x"00",x"00",x"00",x"00",-- 0x38:
   x"00",x"00",x"00",x"00",-- 0x3C:
   x"00",x"00",x"00",x"00",-- 0x40:
   x"00",x"00",x"00",x"00",-- 0x44:
   x"00",x"00",x"00",x"00",-- 0x48:
   x"00",x"00",x"00",x"00",-- 0x4C:
   x"00",x"00",x"00",x"00",-- 0x50:
   x"00",x"00",x"00",x"00",-- 0x54:
   x"00",x"00",x"00",x"00",-- 0x58:
   x"00",x"00",x"00",x"00",-- 0x5C:
   x"00",x"00",x"00",x"00",
   x"00",x"00",x"00",x"00",
   x"00",x"00",x"00",x"00",
   x"00",x"00",x"00",x"00",
   x"00",x"00",x"00",x"00",
   x"00",x"00",x"00",x"00",
   x"00",x"00",x"00",x"00",
   x"00",x"00",x"00",x"00"
   );
begin
process(RAM_CLOCK)
begin
    if(rising_edge(RAM_CLOCK)) then

        if(RAM_WR='1') then -- when write enable = 1,
            -- write input data into RAM at the provided address
            RAM(to_integer(unsigned(RAM_ADDR))) <= RAM_DATA_IN;
            -- The index of the RAM array type needs to be integer so
            -- converts RAM_ADDR from std_logic_vector -> Unsigned -> Interger using numeric_std library
        end if;
    end if;
end process;
 -- Data to be read out
 RAM_DATA_OUT <= RAM(to_integer(unsigned(RAM_ADDR)));
end Behavioral;
